
parameter CTRL_REG_ADDR = 2'b00;
parameter COEFF_REG_ADDR = 2'b01;
parameter SAMPLE_REG_ADDR = 2'b10;
